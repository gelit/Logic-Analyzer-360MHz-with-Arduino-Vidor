
module gla (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
