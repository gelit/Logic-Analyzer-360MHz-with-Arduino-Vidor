
module glb (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
